`default_nettype none

module top (
    input  wire       i_clk,
    input  wire       i_rst,
    output wire [5:0] o_led
);

endmodule
